`ifndef CONTROLSTATES_VH
`define CONTROLSTATES_VH

`define INSTRUCTION_FETCH 4'd0
`define REGISTER_FETCH 4'd1
`define IMMEDIATE_INJECTION3 4'd2
`define ALU_R3 4'd3
`define ALU_RI3 4'd4
`define ALU4 4'd5
`define BRANCH3 4'd6
`define MEMORY_REF3 4'd7
`define LOAD4 4'd8
`define STORE4 4'd9
`define LOAD5 4'd10
`define JUMP3 4'd11

`endif
