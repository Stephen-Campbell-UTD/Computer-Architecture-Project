`timescale 1ns / 1ps
`include "./Control.v"
`include "opcodes.vh"

module testbench ();


  reg [5:0] opcode;
  reg clk;
  wire [3:0] state;

  initial clk <= 0;
  always #5 clk <= ~clk;

  Control uut (
      .opcode(opcode),
      .clk(clk),
      .state(state)
  );

  initial begin
    $dumpfile("./build/main.vcd");
    $dumpvars(0, testbench);
  end


  initial begin
    //ALU R route

    // fist clock ticks at 5ns
    //ALU R takes 4 clocks = 10ns * 4 = 40ns
    // control will be in IF between the beginning of 
    // the 4th clock and end of next clock (35ns to 45ns)
    // IF (0)-> RF (1)-> ALU_R3 (3) -> ALU_4  (5) 
    opcode <= `ADD;
    #40;

    //ALU RI route

    // fist clock ticks at 45ns
    // ALU RI takes 4 clocks = 10ns * 4 = 40ns
    // control will be in IF between the beginning of 
    // the 4th clock and end of next clock (75ns to 85ns)
    // IF (0)-> RF (1)-> ALU_RI3 (4) -> ALU_4  (5) 

    opcode <= `ADDI;
    #40;  //80ns

    //Branch route

    // fist clock ticks at 85ns
    // ALU RI takes 3 clocks = 10ns * 3 = 30ns
    // control will be in IF between the beginning of 
    // the 3th clock and end of next clock (105ns to 115ns)
    // IF (0)-> RF (1)-> BRANCH3 (6)

    opcode <= `BEQ;
    #30;  //110ns

    //Load route

    // fist clock ticks at 115ns
    // Load takes 5 clocks = 10ns * 5 = 50ns
    // control will be in IF between the beginning of 
    // the 5th clock and end of next clock (155ns to 165ns)
    // IF (0)-> RF (1)-> MEMORY_REF3 (7) -> LOAD4 (8) -> LOAD5 (10)

    opcode <= `LD;
    #50;  //160ns

    //Store route

    // fist clock ticks at 165ns
    // Store takes 4 clocks = 10ns * 4 = 40ns
    // control will be in IF between the beginning of 
    // the 4th clock and end of next clock (195ns to 205ns)
    // IF (0)-> RF (1)-> MEMORY_REF3 (7) -> STORE4 (9)
    opcode <= `STR;
    #40;  //200ns

    //Jump route

    // fist clock ticks at 205ns
    // Jump takes 3 clocks = 10ns * 3 = 30ns
    // control will be in IF between the beginning of 
    // the 3rd clock and end of next clock (225ns to 235ns)
    // IF (0)-> RF (1)-> JUMP3 (11)
    opcode <= `JUMP;
    #30;  //230ns

    //Immediate Injection route

    // fist clock ticks at 235ns
    // Imm Injection takes 3 clocks = 10ns * 3 = 30ns
    // control will be in IF between the beginning of 
    // the 3rd clock and end of next clock (265ns to 275ns)
    // IF (0)->  IMMEDIATE_INJECTION3(2)
    opcode <= `LDI;
    #30;  //260ns
    $finish;
  end

endmodule
